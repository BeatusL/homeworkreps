// MY_ISSPE.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module MY_ISSPE (
		input  wire [5:0] probe,      //     probes.probe
		input  wire       source_clk, // source_clk.clk
		output wire [1:0] source      //    sources.source
	);

	altsource_probe_top #(
		.sld_auto_instance_index ("YES"),
		.sld_instance_index      (0),
		.instance_id             ("SP_0"),
		.probe_width             (6),
		.source_width            (2),
		.source_initial_value    ("3"),
		.enable_metastability    ("YES")
	) in_system_sources_probes_0 (
		.source     (source),     //    sources.source
		.source_clk (source_clk), // source_clk.clk
		.probe      (probe),      //     probes.probe
		.source_ena (1'b1)        // (terminated)
	);

endmodule
