
module ISSPE_lab (
	source,
	probe,
	source_clk);	

	output	[1:0]	source;
	input	[3:0]	probe;
	input		source_clk;
endmodule
