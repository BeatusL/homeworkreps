
module SP_unit (
	source,
	probe,
	source_clk);	

	output	[1:0]	source;
	input	[10:0]	probe;
	input		source_clk;
endmodule
