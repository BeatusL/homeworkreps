// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
// Created on Fri Apr 26 00:11:50 2024

// synthesis message_off 10175

`timescale 1ns/1ns

module SM1 (
    clock,reset,x1,x2);

    input clock;
    input reset;
    input x1;
    input x2;
    tri0 reset;
    tri0 x1;
    tri0 x2;
    reg [3:0] fstate;
    reg [3:0] reg_fstate;
    parameter r0=0,r1=1,r2=2,r3=3;

    always @(posedge clock or negedge reset)
    begin
        if (~reset) begin
            fstate <= r0;
        end
        else begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or x1 or x2)
    begin
        case (fstate)
            r0: begin
                if ((~(x2) & ~(x1)))
                    reg_fstate <= r2;
                else if ((~(x2) & x1))
                    reg_fstate <= r1;
                else if ((x2 & x1))
                    reg_fstate <= r3;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= r0;
            end
            r1: begin
                if ((~(x2) & ~(x1)))
                    reg_fstate <= r2;
                else if ((x2 & x1))
                    reg_fstate <= r3;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= r1;
            end
            r2: begin
                if ((~(x2) & ~(x1)))
                    reg_fstate <= r2;
                else if ((~(x2) & x1))
                    reg_fstate <= r1;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= r2;
            end
            r3: begin
                if ((~(x2) & ~(x1)))
                    reg_fstate <= r1;
                else if ((x2 & x1))
                    reg_fstate <= r0;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= r3;
            end
            default: begin
                $display ("Reach undefined state");
            end
        endcase
    end
endmodule // SM1
