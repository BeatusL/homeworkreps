-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Fri Apr 05 21:46:45 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SM1 IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        x1 : IN STD_LOGIC := '0';
        x2 : IN STD_LOGIC := '0'
    );
END SM1;

ARCHITECTURE BEHAVIOR OF SM1 IS
    TYPE type_fstate IS (r0,r1,r2,r3);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='0') THEN
            fstate <= r0;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,x1,x2)
    BEGIN
        CASE fstate IS
            WHEN r0 =>
                IF ((NOT((x2 = '1')) AND NOT((x1 = '1')))) THEN
                    reg_fstate <= r2;
                ELSIF ((NOT((x2 = '1')) AND (x1 = '1'))) THEN
                    reg_fstate <= r1;
                ELSIF (((x2 = '1') AND (x1 = '1'))) THEN
                    reg_fstate <= r3;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= r0;
                END IF;
            WHEN r1 =>
                IF ((NOT((x2 = '1')) AND NOT((x1 = '1')))) THEN
                    reg_fstate <= r2;
                ELSIF (((x2 = '1') AND (x1 = '1'))) THEN
                    reg_fstate <= r3;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= r1;
                END IF;
            WHEN r2 =>
                IF ((NOT((x2 = '1')) AND NOT((x1 = '1')))) THEN
                    reg_fstate <= r2;
                ELSIF ((NOT((x2 = '1')) AND (x1 = '1'))) THEN
                    reg_fstate <= r1;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= r2;
                END IF;
            WHEN r3 =>
                IF ((NOT((x2 = '1')) AND NOT((x1 = '1')))) THEN
                    reg_fstate <= r1;
                ELSIF (((x2 = '1') AND (x1 = '1'))) THEN
                    reg_fstate <= r0;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= r3;
                END IF;
            WHEN OTHERS => 
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
